//---------------------------Galileo University---------------------------//
//	Main Collaborators:
//	- Rodrigo Cordero
//	- Kevin Hernandez
//
//	Module Name: riscv.v
//	Project: FPGA RISC V
//	Description: Verilog module which describes the behavior of a RISC V processor
//
//
//	Update History:
//	- 01/14/2019: Creation of the module
//
//-------------------------------------------------------------------------//

module riscv(clk, fetch_addr, instruction, result);
	input clk;
	output [31:0] fetch_addr, instruction, result;

	

endmodule