module and32bits(A,B,C);
  input [31:0] A,B;
  output [31:0] C;
  	//Spam de ANDs
	and(C[0], A[0], B[0]);
	and(C[1], A[1], B[1]);
	and(C[2], A[2], B[2]);
	and(C[3], A[3], B[3]);
	and(C[4], A[4], B[4]);
	and(C[5], A[5], B[5]);
	and(C[6], A[6], B[6]);
	and(C[7], A[7], B[7]);
	and(C[8], A[8], B[8]);
	and(C[9], A[9], B[9]);
	and(C[10], A[10], B[10]);
	and(C[11], A[11], B[11]);
	and(C[12], A[12], B[12]);
	and(C[13], A[13], B[13]);
	and(C[14], A[14], B[14]);
	and(C[15], A[15], B[15]);
	and(C[16], A[16], B[16]);
	and(C[17], A[17], B[17]);
	and(C[18], A[18], B[18]);
	and(C[19], A[19], B[19]);
	and(C[20], A[20], B[20]);
	and(C[21], A[21], B[21]);
	and(C[22], A[22], B[22]);
	and(C[23], A[23], B[23]);
	and(C[24], A[24], B[24]);
	and(C[25], A[25], B[25]);
	and(C[26], A[26], B[26]);
	and(C[27], A[27], B[27]);
	and(C[28], A[28], B[28]);
	and(C[29], A[29], B[29]);
	and(C[30], A[30], B[30]);
	and(C[31], A[31], B[31]);
endmodule

module or32bits(A,B,C);
  input [31:0] A,B;
  output [31:0] C;
  	//Spam de ORs
	or(C[0], A[0], B[0]);
	or(C[1], A[1], B[1]);
	or(C[2], A[2], B[2]);
	or(C[3], A[3], B[3]);
	or(C[4], A[4], B[4]);
	or(C[5], A[5], B[5]);
	or(C[6], A[6], B[6]);
	or(C[7], A[7], B[7]);
	or(C[8], A[8], B[8]);
	or(C[9], A[9], B[9]);
	or(C[10], A[10], B[10]);
	or(C[11], A[11], B[11]);
	or(C[12], A[12], B[12]);
	or(C[13], A[13], B[13]);
	or(C[14], A[14], B[14]);
	or(C[15], A[15], B[15]);
	or(C[16], A[16], B[16]);
	or(C[17], A[17], B[17]);
	or(C[18], A[18], B[18]);
	or(C[19], A[19], B[19]);
	or(C[20], A[20], B[20]);
	or(C[21], A[21], B[21]);
	or(C[22], A[22], B[22]);
	or(C[23], A[23], B[23]);
	or(C[24], A[24], B[24]);
	or(C[25], A[25], B[25]);
	or(C[26], A[26], B[26]);
	or(C[27], A[27], B[27]);
	or(C[28], A[28], B[28]);
	or(C[29], A[29], B[29]);
	or(C[30], A[30], B[30]);
	or(C[31], A[31], B[31]);
endmodule

module xor32bits(A,B,C);
  input [31:0] A,B;
  output [31:0] C;
  	//Spam de XORs
	xor(C[0], A[0], B[0]);
	xor(C[1], A[1], B[1]);
	xor(C[2], A[2], B[2]);
	xor(C[3], A[3], B[3]);
	xor(C[4], A[4], B[4]);
	xor(C[5], A[5], B[5]);
	xor(C[6], A[6], B[6]);
	xor(C[7], A[7], B[7]);
	xor(C[8], A[8], B[8]);
	xor(C[9], A[9], B[9]);
	xor(C[10], A[10], B[10]);
	xor(C[11], A[11], B[11]);
	xor(C[12], A[12], B[12]);
	xor(C[13], A[13], B[13]);
	xor(C[14], A[14], B[14]);
	xor(C[15], A[15], B[15]);
	xor(C[16], A[16], B[16]);
	xor(C[17], A[17], B[17]);
	xor(C[18], A[18], B[18]);
	xor(C[19], A[19], B[19]);
	xor(C[20], A[20], B[20]);
	xor(C[21], A[21], B[21]);
	xor(C[22], A[22], B[22]);
	xor(C[23], A[23], B[23]);
	xor(C[24], A[24], B[24]);
	xor(C[25], A[25], B[25]);
	xor(C[26], A[26], B[26]);
	xor(C[27], A[27], B[27]);
	xor(C[28], A[28], B[28]);
	xor(C[29], A[29], B[29]);
	xor(C[30], A[30], B[30]);
	xor(C[31], A[31], B[31]);
endmodule
