//---------------------------Galileo University---------------------------//
//	Main Collaborators:
//	- Rodrigo Cordero
//	- Kevin Hernandez
//
//	Module Name: controll.v
//	Project: FPGA RISC V
//	Description: Verilog module which describes the behaviour for Risc V's Controll section.
//
//
//	Update History:
//	- 02/01/2019: Creation of the module and the following submodules: immGenSelector, muxABSelector,
//								writeRegEnable, loadEnable, writeBack and pcEnable
//	- 03/01/2019: Added a submodule description and the following submodules: unsignedOperations
//
//	-04/01/2019: Added LoadControll, AluSelector, BranchSelector submodules and their connections. Also added the 2nd stage of the pipeline

//
//	Submodule Description:
//	- immGenSelector:	The purpose of this submodule is to send a signal to the Immediate Generator 
//
//-------------------------------------------------------------------------//

module controll(clk, instruction, );
	input clk, blt, beq;
	input [31:0] instruction;
	//*************
	output reg [3:0] ALUSelector;
	output reg BrUnsigned, Bres, nop, WMemEnable;
	output reg [1:0] LoadSelector;
	reg [3:0] wALUSelector;
	reg wNop = 1'b0;
	reg wandor, Inst6, Inst2, WME1;
	reg [31:0] wBControll;
	reg [1:0] wLoadS, loadControll;
	ALUSel aS(instruction, wALUSelector);
	loadControll lC(instruction, loadControll);
	brControll BC1(wBControll, blt, beq, Bres);
	//**********

	reg pipelines [0:7];
	always @ (posedge clk)
	fork
		//-----Immediate Generator Selector-----//
		begin
			//*****
			ALUSelector = wALUSelector;
			BrUnsigned = instruction[13];
			if(~wNop)
				begin
					wBControll = instruction;
					wandor = ((instruction[6] & instruction[2]) | (Bres & instruction[6] & ~instruction[2]));
				end
			else if(wNop)
				begin
					wandor = 1'b0;
					wBControll = 32'b0;
					WME1 = 1'b0;
				end
			nop = wandor;
			wNop = wandor;
			LoadSelector = wLoadS;
			wLoadS = loadControll;
			WMemEnable = WME1;
			WME1 = WME;
			//*****
		end


	join
endmodule

module immGenSelector(clk, nop, opcode, pipeline);
	//-----Immediate Generator Selector-----//
	input clk, nop;
	input [6:0] opcode;
	output [4:0] pipeline;

	reg [4:0] pipeline;

	always @ (posedge clk)
		if(nop)
			fork
				pipeline[0] = 0;																		//Type I
				pipeline[1] = 0;																		//Type S
				pipeline[2] = 0;																		//Type U
				pipeline[3] = 0;																		//Type SB
				pipeline[4] = 0;																		//Type UJ
			join
		else
			fork
				pipeline[0] = (~opcode[5] & ~opcode[2]) | (~opcode[4] & ~opcode[3] & opcode[2]);							//Type I
				pipeline[1] = ~opcode[6] & opcode[5] & ~opcode[4];	//Type S
				pipeline[2] = ~opcode[6] & opcode[2];								//Type U
				pipeline[3] = opcode[6] & ~opcode[3] & ~opcode[2];	//Type SB
				pipeline[4] = opcode[3];														//Type UJ
			join
endmodule

module muxABSelector(clk, nop, opcode, pipeline);
	//-----Selector for multiplexor A and B-----//
	input clk, nop;
	input [6:0] opcode;
	output [1:0] pipeline;

	reg [1:0] pipeline;

	always @ (posedge clk)
		if(nop)
			fork
				pipeline[0] = 0;																																				//Multiplexor A
				pipeline[1] = 0;																																				//Multiplexor B
			join
		else
			fork
				pipeline[0] = ~((~opcode[6] & ~opcode[2]) | (~opcode[4] & ~opcode[3] & opcode[2]));			//Multiplexor A
				pipeline[1] = ~(opcode[5] & opcode[4] & ~opcode[2]);																		//Multiplexor B
			join
endmodule

module writeRegEnable(clk, nop, opcode, pipeline3);
	//-----Write Register Enable signal-----//
	input clk, nop;
	input [6:0] opcode;
	output pipeline3;

	reg pipeline, pipeline2, pipeline3;

	always @ (posedge clk)
	begin
		pipeline3 = pipeline2;
		pipeline2 = pipeline;
		if(nop)
			pipeline = 0;
		else
			pipeline = (~opcode[5] | opcode[4] | opcode[2]) & opcode[1] & opcode[0];
	end
endmodule

module writeMemEnable(clk, nop, opcode, pipeline2);
	//-----Write Memory Enable signal-----//
	input clk, nop;
	input [6:0] opcode;
	output pipeline2;

	reg pipeline, pipeline2;

	always @ (posedge clk)
	begin
		pipeline2 = pipeline;
		if(nop)
			pipeline = 0;
		else
			pipeline = ~opcode[6] & opcode[5] & ~opcode[4];
	end
endmodule

module loadEnable(clk, opcode, pipeline2);
	//-----Load Enable signal-----//
	input clk;
	input [6:0] opcode;
	output pipeline2;

	reg pipeline, pipeline2;

	always @ (posedge clk)
	begin
		pipeline2 = pipeline;
		pipeline = ~opcode[6] & ~opcode[5] & ~opcode[4] & ~opcode[3] & ~opcode[2] & opcode[1] & opcode[0];
    end
endmodule

module writeBack(clk, opcode, pipeline2);
	//-----Write Back signal-----//
	input clk;
	input [6:0] opcode;
	output [1:0] pipeline2;

	reg [1:0] pipeline, pipeline2;

	always @ (posedge clk)
	begin
		pipeline2 = pipeline;
		if(~opcode[6] & opcode[5] & opcode[2])
			pipeline = 2'b11;
		else if(~opcode[5] & ~opcode[4])
			pipeline = 2'b10;
		else if((opcode[4] & ~opcode[2]) | (~opcode[5] & opcode[2]))
			pipeline = 2'b01;
		else
			pipeline = 2'b00;
	end
endmodule

module pcEnable(clk, nop, bres, opcode, pipeline2);
	//-----PC Enable signal-----//
	input clk, nop, bres;
	input [6:0] opcode;
	output pipeline2;

	reg [6:0] pipeline;
	reg pipeline2;

	always @ (posedge clk)
	begin
		pipeline2 = (bres | pipeline[2]) & pipeline[6];
		if(nop)
			pipeline = 7'b0000000;
		else
			pipeline = opcode;
	end
endmodule

module unsignedOperations(clk, nop, instruction);
	//-----Unsigned Operations for ALU signal-----//
	input clk, nop;
	input [31:0] instruction;
	output pipeline;

	reg pipeline;

	always @ (posedge clk)
	if(nop)
		pipeline = 0;
	else
		pipeline = ((~instruction[30] & instruction[14] & ~instruction[13]) | (~instruction[14] & instruction[13])) & instruction[12] & instruction[4] & ~instruction[2];
endmodule

module loadControll(input [31:0] Inst,
                    output reg [1:0] loadMux);
  
  always @(Inst)
    case ({Inst[14], Inst[13], Inst[12]})
      3'b000: loadMux = 0;
      3'b001: loadMux = 1;
      3'b010: loadMux = 2;
      default: loadMux = 0;
    endcase
endmodule

module ALUSel(input [31:0] Inst,
              output reg [3:0] ALUSelOut);
  
  reg wiSll, wiSlr, wiAdd, wiAnd1, wiAnd2, wiAnd3, wiAnd4, wiOr, wiXor, wiMul, wiMulh, wiDiv, wiRem, wiSub, wiSlt;
  
  always @(Inst)
      fork
        case (Inst[0] & Inst[1])
          1'b0 : ALUSelOut = 2;
          1'b1 : 
            begin
              wiSll = 1'b0; //Sll
              
              wiSlr = Inst[14] & ~Inst[13] & Inst[12] & Inst[4] & ~Inst[2]; // Slr
            
              wiAdd = (((~Inst[14] & ~Inst[13] & ~Inst[12] & Inst[4]) & ((~Inst[30] & ~Inst[25] & Inst[5] & ~Inst[2]) |  ~Inst[5])) | ~Inst[4]);
            
              wiAnd1 = (Inst[14] & Inst[13] & Inst[12] & Inst[4]);
              wiAnd2 = (Inst[5] & ~Inst[2]);
              wiAnd3 = wiAnd1 | wiAnd2;
              wiAnd4 = wiAnd1 & wiAnd3; //And
            
               wiOr = ((Inst[14] & Inst[13] & ~Inst[12] & Inst[4] & ((~Inst[25] & Inst[5] & ~Inst[2]) | ~Inst[5]))); // Or
            
               wiXor = ((Inst[14] & ~Inst[13] & ~Inst[12] & Inst[4] & ((~Inst[25] & Inst[5] & ~Inst[2]) | ~Inst[5]))); // Xor
            
              wiSlt = (~Inst[14] & Inst[13] & Inst[4] & ~Inst[2]); // Slt
            
              wiMul = ((~Inst[14] & ~Inst[13] & ~Inst[12] & Inst[4] & ~Inst[30] & Inst[25] & Inst[5] & ~Inst[2])); // Mul
            
              wiMulh = (~Inst[14] & ~Inst[13] & Inst[12] & Inst[4] & Inst[25] & Inst[5] & ~Inst[2]); // Mulh
            
              wiDiv = ((Inst[14] & ~Inst[13] & ~Inst[12] & Inst[4] & Inst[25] & Inst[5] & ~Inst[2])); // Div
            
              wiRem = ((Inst[14] & Inst[13] & ~Inst[12] & Inst[4] & Inst[25] & Inst[5] & ~Inst[2])); // Rem
            
              wiSub = ((~Inst[14] & ~Inst[13] & ~Inst[12] & Inst[4] & Inst[30] & ~Inst[25] & Inst[5] & ~Inst[2])); // Sub
              
              
              ALUSelOut = wiSll | (wiSlr * 1) | (wiAdd * 2) | (wiAnd4 * 3) | (wiOr * 4) | (wiXor * 5) | (wiMul * 7) |  (wiMulh * 8) | (wiDiv * 9) | (wiRem * 10) | (wiSub * 11) | (wiSlt * 6);
            end
        endcase
      join
endmodule

module brControll(input [31:0] Inst,
                  input blt, beq, 
                  output reg result);
  
  always @(Inst)
      fork
        case(~Inst[12])
          1'b0:
            begin
              if(~Inst[14])
                result = ~beq;
              else
                result = ~blt;
            end
          1'b1:
              begin
                if(~Inst[14])
                  result = beq;
                else
                  result = blt;
              end
        endcase
      join
                
endmodule
