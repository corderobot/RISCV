module ShiftLogico12BitIzquierda(Original, Nuevo);
  input [31:0] Original;
  output [31:0] Nuevo;
  and (Nuevo[0], 1'b0, 1'b1);
  and (Nuevo[1], 1'b0, 1'b1);
  and (Nuevo[2], 1'b0, 1'b1);
  and (Nuevo[3], 1'b0, 1'b1);
  and (Nuevo[4], 1'b0, 1'b1);
  and (Nuevo[5], 1'b0, 1'b1);
  and (Nuevo[6], 1'b0, 1'b1);
  and (Nuevo[7], 1'b0, 1'b1);
  and (Nuevo[8], 1'b0, 1'b1);
  and (Nuevo[9], 1'b0, 1'b1);
  and (Nuevo[10], 1'b0, 1'b1);
  and (Nuevo[11], 1'b0, 1'b1);
  and (Nuevo[12], Original[0], 1'b1);
  and (Nuevo[13], Original[1], 1'b1);
  and (Nuevo[14], Original[2], 1'b1);
  and (Nuevo[15], Original[3], 1'b1);
  and (Nuevo[16], Original[4], 1'b1);
  and (Nuevo[17], Original[5], 1'b1);
  and (Nuevo[18], Original[6], 1'b1);
  and (Nuevo[19], Original[7], 1'b1);
  and (Nuevo[20], Original[8], 1'b1);
  and (Nuevo[21], Original[9], 1'b1);
  and (Nuevo[22], Original[10], 1'b1);
  and (Nuevo[23], Original[11], 1'b1);
  and (Nuevo[24], Original[12], 1'b1);
  and (Nuevo[25], Original[13], 1'b1);
  and (Nuevo[26], Original[14], 1'b1);
  and (Nuevo[27], Original[15], 1'b1);
  and (Nuevo[28], Original[16], 1'b1);
  and (Nuevo[29], Original[17], 1'b1);
  and (Nuevo[30], Original[18], 1'b1);
  and (Nuevo[31], Original[19], 1'b1);
endmodule;
