// Módulos
